///////////////////////////////////////////////////////////////////////////////
// File: power_control.sv
// Date: 2026.02.03
// Designer: drake.lee
// Description: Power control module for ROIC bias voltage sequencing
//              Extracted from cyan_top.sv (Week 8 - M8-2)
//
// Functionality:
//   - Power sequencing control for ROIC initialization
//   - Bias voltage control (VBIAS, AVDD1, AVDD2)
//   - Power-on initialization coordination with init module
//   - Reset generation for power control FSM
//
// Revision History:
//    2026.02.04 - RST-004 fix: Removed incorrect init_rst output (generated by init module)
//    2026.02.03 - Initial extraction from cyan_top.sv
//
///////////////////////////////////////////////////////////////////////////////

module power_control (
    // Clock and Reset
    input  logic        clk_20mhz,
    input  logic        rst_n_20mhz,          // Active-LOW reset

    // Power Initialization Control (from init module)
    input  logic        pwr_init_step1,       // Power init step 1 enable
    input  logic        pwr_init_step2,       // Power init step 2 enable
    input  logic        pwr_init_step3,       // Power init step 3 enable
    input  logic        pwr_init_step4,       // Power init step 4 enable
    input  logic        pwr_init_step5,       // Power init step 5 enable
    input  logic        pwr_init_step6,       // Power init step 6 enable

    // Back Bias Control (from roic_gate_drv_gemini)
    input  logic        back_bias,            // Back bias signal from gate driver

    // FSM Reset Control
    output logic        fsm_rst_index,        // FSM reset index output

    // ROIC Bias Power Outputs
    output logic        ROIC_VBIAS,           // ROIC bias voltage output
    output logic        ROIC_AVDD1,           // ROIC AVDD1 power output
    output logic        ROIC_AVDD2            // ROIC AVDD2 power output
);

    //==========================================================================
    // Internal Signals
    //==========================================================================
    logic fsm_drv_rst;              // FSM driver reset (active-LOW)

    //==========================================================================
    // FSM Reset Generation
    //==========================================================================
    // FSM driver reset is active-LOW, controlled by rst_n_20mhz and FSM reset index
    assign fsm_drv_rst = rst_n_20mhz & ~fsm_rst_index;

    // Note: init_rst is generated by the init module, not power_control
    // RST-004 fix: Removed incorrect init_rst output from this module

    //==========================================================================
    // Power Sequencing Control
    //==========================================================================
    // The power sequencing follows these steps during initialization:
    // Step 1: Enable ROIC_AVDD1 (first power rail)
    // Step 2: Enable ROIC_AVDD2 (second power rail)
    // Step 3-6: Additional power sequencing steps (internal to init module)
    //
    // The power rails are enabled when:
    //   1. The corresponding init step is active
    //   2. Power down is not asserted
    //
    // Power rail outputs:
    assign ROIC_AVDD1 = pwr_init_step1;
    assign ROIC_AVDD2 = pwr_init_step2;

    //==========================================================================
    // Bias Voltage Control
    //==========================================================================
    // ROIC_VBIAS is controlled by the back_bias signal from the gate driver.
    // This signal is generated by roic_gate_drv_gemini based on the
    // back_bias FSM state and controls the bias voltage applied to the ROIC.
    assign ROIC_VBIAS = back_bias;

    //==========================================================================
    // Notes on Power Sequencing
    //==========================================================================
    // Power-on sequence (controlled by init module):
    //   1. pwr_init_step1 -> Enables AVDD1
    //   2. pwr_init_step2 -> Enables AVDD2
    //   3. pwr_init_step3-6 -> Internal sequencing steps
    //
    // Power-off sequence (reverse order):
    //   1. Step 6 -> 3 disabled
    //   2. pwr_init_step2 disabled -> AVDD2 off
    //   3. pwr_init_step1 disabled -> AVDD1 off
    //
    // The back_bias signal is controlled independently by the gate driver
    // based on the FSM back_bias_index state.

endmodule
